//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.01 (64-bit)
//Part Number: GW5A-LV25UG324ES
//Device: GW5A-25
//Device Version: A
//Created Time: Sun Sep 22 20:16:25 2024

module fft_rom1 (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0A7607BF089B0BAC0C8409C6070607D90AE10BB208ED062806F609FA0AC70800;
defparam prom_inst_0.INIT_RAM_01 = 256'h0DA60B1A088B098D0CC30DC00B260889097E0CA70D960AEE0844092C0C470D2A;
defparam prom_inst_0.INIT_RAM_02 = 256'h0AE70C0B099A072808490B9F0CBE0A4707CE08E80C370D4D0ACC084909590C9C;
defparam prom_inst_0.INIT_RAM_03 = 256'h057708C509DF076704F0060F09650A87081505A406C70A220B4708D70668078D;
defparam prom_inst_0.INIT_RAM_04 = 256'h04120502082A0920068303EA04E7081E09210692040605100854096306E10461;
defparam prom_inst_0.INIT_RAM_05 = 256'h08B005ED06BE09C70A9B07DC051E05F7090809E4072F047B055F087A096306B9;
defparam prom_inst_0.INIT_RAM_06 = 256'h0E130B560898096C0C750D460A8307BE088D0B920C60099A06D307A20AA60B75;
defparam prom_inst_0.INIT_RAM_07 = 256'h0E410F3F0CA60A0B0B010E2A0F1B0C7409CB0AB40DD00EB40C01094C0A290D3A;
defparam prom_inst_0.INIT_RAM_08 = 256'h09B00D080E280BB3093C0A570DA70EBE0C3F09BE0ACE0E130F1E0C930A050B09;
defparam prom_inst_0.INIT_RAM_09 = 256'h063E075E0AB60BD9096906FA081F0B7B0CA20A3407C608EC0C490D6E0AFE088E;
defparam prom_inst_0.INIT_RAM_0A = 256'h07B4051C061C09540A5907CC0542064E09930AA5082405A606BE0A0E0B2A08B3;
defparam prom_inst_0.INIT_RAM_0B = 256'h0BAB08EE0633070E0A210AFF084C059A0680099D0A8707E0053B062C09570A4E;
defparam prom_inst_0.INIT_RAM_0C = 256'h0D620E360B7508B309840C8B0D5B0A9707D308A30BAA0C7B09B806F707CA0AD5;
defparam prom_inst_0.INIT_RAM_0D = 256'h0BC90EF50FE80D440A9D0B880EA70F8D0CDC0A2A0B090E1C0EF80C3D09810A57;
defparam prom_inst_0.INIT_RAM_0E = 256'h09DD0AFB0E4D0F670CEA0A6B0B7E0EC50FD30D4B0ABF0BC60EFF10000D6A0AD1;
defparam prom_inst_0.INIT_RAM_0F = 256'h09E10775089D0BFB0D240AB9084E09770CD50DFD0B9009220A480DA20EC50C52;
defparam prom_inst_0.INIT_RAM_10 = 256'h0AA7081D059506A409EC0B000882060607210A740B92091E06AB07CF0B290C4F;
defparam prom_inst_0.INIT_RAM_11 = 256'h0A440B25087405C606AE09CE0ABB08160573066809950A8F07F705620664099F;
defparam prom_inst_0.INIT_RAM_12 = 256'h097C0C850D580A9707D608A90BB20C8609C6070707DD0AEB0BC409090651072E;
defparam prom_inst_0.INIT_RAM_13 = 256'h0A6A0B570E790F620CB40A040AE60DFC0EDA0C2209680A410D4F0E260B6708A8;
defparam prom_inst_0.INIT_RAM_14 = 256'h0C8C0A100B260E6F0F800CFA0A710B7A0EB70FBA0D260A900B8B0EBA0FAF0D0E;
defparam prom_inst_0.INIT_RAM_15 = 256'h0C9D0A3407CB08F70C580D830B1808AD09D50D310E570BE609740A950DEA0F06;
defparam prom_inst_0.INIT_RAM_16 = 256'h093C0A5207D7055E067B09D00AF1087F060F07350A920BBB094F06E508100B71;
defparam prom_inst_0.INIT_RAM_17 = 256'h05D708FA09E9074604A6059D08CD09C9073404A105A608E309ED076504E005F2;
defparam prom_inst_0.INIT_RAM_18 = 256'h06DB07B00ABB0B9108D4061706F00A000ADA0823056C064C09640A48079904ED;
defparam prom_inst_0.INIT_RAM_19 = 256'h0B9708E909CD0CE50DC50B0F085809330C430D1C0A5F07A208780B840C59099A;
defparam prom_inst_0.INIT_RAM_1A = 256'h0E440BC009390A440D820E870BF609610A5E0D8F0E860BE709450A350D580E43;
defparam prom_inst_0.INIT_RAM_1B = 256'h0B000C2C09C4075A08830BE20D090A9A082A094C0CA30DC10B4908CE09E60D31;
defparam prom_inst_0.INIT_RAM_1C = 256'h050B08610984071404A505CC092B0A5507EB058206AE0A110B3E08D70670079D;
defparam prom_inst_0.INIT_RAM_1D = 256'h0321041A074B084805B4032304280767087205EC0368047B07C608DE066403EC;
defparam prom_inst_0.INIT_RAM_1E = 256'h073E0483055C086D0949069203DD04BE07D608BB060E0362044E0772086205C0;
defparam prom_inst_0.INIT_RAM_1F = 256'h0C23096E06B707930AA40B7D08C2060506DC09E80ABE080005420618092409FB;
defparam prom_inst_0.INIT_RAM_20 = 256'h0BD80CDD0A4C07B808B50BE60CDF0A40079E088E0BB20C9E09F20745082A0B42;
defparam prom_inst_0.INIT_RAM_21 = 256'h06D50A340B5B08EC067C079F0AF50C14099C0722083A0B850C980A14078E0899;
defparam prom_inst_0.INIT_RAM_22 = 256'h02F7041E077D08A6063C03D4050008630990072904C205EF09520A7E081505AB;
defparam prom_inst_0.INIT_RAM_23 = 256'h040A0179027E05BC06C7044001BC02CF061A073204B7023F035D06B407D60566;
defparam prom_inst_0.INIT_RAM_24 = 256'h07A804F1023B031B06330717046901BD02A805CB06BB0419017A027105A2069F;
defparam prom_inst_0.INIT_RAM_25 = 256'h091009E9072C046F054508500925066603A7047C0788085E05A102E403BD06CD;
defparam prom_inst_0.INIT_RAM_26 = 256'h07330A630B5A08BA061707060A290B13086705B8069C09B40A9407DD05260600;
defparam prom_inst_0.INIT_RAM_27 = 256'h050F063009850AA2082905AE06C40A0E0B20089B0613071D0A5A0B5F08CC0637;
defparam prom_inst_0.INIT_RAM_28 = 256'h04E8027D03A80709083505CC0363048F07F0091B06B10445056E08CB09F10781;
defparam prom_inst_0.INIT_RAM_29 = 256'h058F03060080019104DA05F0037400FA0216056B068C041A01A902CF062B0753;
defparam prom_inst_0.INIT_RAM_2A = 256'h051A05FC034C009E018704A9059602F2005101460475057002DA004601490486;
defparam prom_inst_0.INIT_RAM_2B = 256'h044E0757082A056902A8037B06840758049901DA02B105BF069803DE01260204;
defparam prom_inst_0.INIT_RAM_2C = 256'h0545063209520A3A078C04DB05BC08D209AF06F7043C0515082308F9063A037A;
defparam prom_inst_0.INIT_RAM_2D = 256'h077E05000614095C0A6B07E305590661099C0A9E08090571066B09980A8D07EA;
defparam prom_inst_0.INIT_RAM_2E = 256'h07B2054702DC04050763088B061F03B104D70831095506E2046E058C08DF09FA;
defparam prom_inst_0.INIT_RAM_2F = 256'h048205950316009901B30505062303AE013B025E05B806DE04700203032B0689;
defparam prom_inst_0.INIT_RAM_30 = 256'h01590478056302BC0018010B0437052F029600000101043A054102B5002D013B;
defparam prom_inst_0.INIT_RAM_31 = 256'h02A50375067C074D048B01CA029E05A9067F03C3010801E404F705D603240073;
defparam prom_inst_0.INIT_RAM_32 = 256'h07B4050105DF08F209CD07120455052B08360909064803850456075D082D0569;
defparam prom_inst_0.INIT_RAM_33 = 256'h0ABE083405A706AC09E40AE4084C05B206A909D40AC508200579066309800A66;
defparam prom_inst_0.INIT_RAM_34 = 256'h07E1090606970427054A08A209C2074D04D605F209420A5A07DC055B066D09B2;
defparam prom_inst_0.INIT_RAM_35 = 256'h025905A906C4044D01D802F8065007720502029203B70714083A05CC035E0485;
defparam prom_inst_0.INIT_RAM_36 = 256'h00E501D604FF05F5035A00C101BF04F705FB036D00E201ED0532064203C10142;
defparam prom_inst_0.INIT_RAM_37 = 256'h057D02BA038B0694076804AA01ED02C605D706B403FF014C0230054C0635038C;
defparam prom_inst_0.INIT_RAM_38 = 256'h0AE208240565063909420A130750048B055A085E092D066603A0046E07730842;
defparam prom_inst_0.INIT_RAM_39 = 256'h0B190C16097D06E007D60AFE0BEE0947069D07860AA10B8508D1061C06F80A09;
defparam prom_inst_0.INIT_RAM_3A = 256'h069B09F10B1008990621073B0A890B9F091F069D07AC0AF00BFA096E06DF07E2;
defparam prom_inst_0.INIT_RAM_3B = 256'h0342046107B708D8066603F5051908730998072904B905DE09390A5C07EB0579;
defparam prom_inst_0.INIT_RAM_3C = 256'h04DA0240033D0673077504E6025A036406A707B7053402B303C90718083205B9;
defparam prom_inst_0.INIT_RAM_3D = 256'h08FA063A037C045407650841058A02D603B906D407BC0512026A035906820777;
defparam prom_inst_0.INIT_RAM_3E = 256'h0AE10BB208ED062806F609FA0AC7080005390606090A09D80713044E051F0827;
defparam prom_inst_0.INIT_RAM_3F = 256'h097E0CA70D960AEE0844092C0C470D2A0A7607BF089B0BAC0C8409C6070607D9;

endmodule //fft_rom1
