//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.01 (64-bit)
//Part Number: GW5A-LV25UG324ES
//Device: GW5A-25
//Device Version: A
//Created Time: Fri Sep 20 18:14:50 2024

module fft_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0A91094B0B770F0E0EE809DD04D104A508330A5208FB07A309BF0D480D150800;
defparam prom_inst_0.INIT_RAM_01 = 256'h0FD50B050631063C09FF0C520B2C0A040C4D10000FF50B05061105FD09A10BD5;
defparam prom_inst_0.INIT_RAM_02 = 256'h077109F108FB08040A810E690E9509DD0524054A09290B990A9109870BEF0FC1;
defparam prom_inst_0.INIT_RAM_03 = 256'h06D70AB60ADC0623016B0197057F07FC0705060F088F0C7C0CAF080003510384;
defparam prom_inst_0.INIT_RAM_04 = 256'h000B000003B305FC04D403AE060109C409CF04FB002B003F04110679056F0467;
defparam prom_inst_0.INIT_RAM_05 = 256'h070505AE07CD0B5B0B2F0623011800F2048906B5056F042B065F0A0309EF04FB;
defparam prom_inst_0.INIT_RAM_06 = 256'h0EE809DD04D104A508330A5208FB07A309BF0D480D15080002EB02B80641085D;
defparam prom_inst_0.INIT_RAM_07 = 256'h09FF0C520B2C0A040C4D10000FF50B05061105FD09A10BD50A91094B0B770F0E;
defparam prom_inst_0.INIT_RAM_08 = 256'h0A810E690E9509DD0524054A09290B990A9109870BEF0FC10FD50B050631063C;
defparam prom_inst_0.INIT_RAM_09 = 256'h016B0197057F07FC0705060F088F0C7C0CAF080003510384077109F108FB0804;
defparam prom_inst_0.INIT_RAM_0A = 256'h04D403AE060109C409CF04FB002B003F04110679056F046706D70AB60ADC0623;
defparam prom_inst_0.INIT_RAM_0B = 256'h0B2F0623011800F2048906B5056F042B065F0A0309EF04FB000B000003B305FC;
defparam prom_inst_0.INIT_RAM_0C = 256'h08330A5208FB07A309BF0D480D15080002EB02B80641085D070505AE07CD0B5B;
defparam prom_inst_0.INIT_RAM_0D = 256'h0C4D10000FF50B05061105FD09A10BD50A91094B0B770F0E0EE809DD04D104A5;
defparam prom_inst_0.INIT_RAM_0E = 256'h0524054A09290B990A9109870BEF0FC10FD50B050631063C09FF0C520B2C0A04;
defparam prom_inst_0.INIT_RAM_0F = 256'h0705060F088F0C7C0CAF080003510384077109F108FB08040A810E690E9509DD;
defparam prom_inst_0.INIT_RAM_10 = 256'h09CF04FB002B003F04110679056F046706D70AB60ADC0623016B0197057F07FC;
defparam prom_inst_0.INIT_RAM_11 = 256'h048906B5056F042B065F0A0309EF04FB000B000003B305FC04D403AE060109C4;
defparam prom_inst_0.INIT_RAM_12 = 256'h09BF0D480D15080002EB02B80641085D070505AE07CD0B5B0B2F0623011800F2;
defparam prom_inst_0.INIT_RAM_13 = 256'h061105FD09A10BD50A91094B0B770F0E0EE809DD04D104A508330A5208FB07A3;
defparam prom_inst_0.INIT_RAM_14 = 256'h0A9109870BEF0FC10FD50B050631063C09FF0C520B2C0A040C4D10000FF50B05;
defparam prom_inst_0.INIT_RAM_15 = 256'h0CAF080003510384077109F108FB08040A810E690E9509DD0524054A09290B99;
defparam prom_inst_0.INIT_RAM_16 = 256'h04110679056F046706D70AB60ADC0623016B0197057F07FC0705060F088F0C7C;
defparam prom_inst_0.INIT_RAM_17 = 256'h065F0A0309EF04FB000B000003B305FC04D403AE060109C409CF04FB002B003F;
defparam prom_inst_0.INIT_RAM_18 = 256'h02EB02B80641085D070505AE07CD0B5B0B2F0623011800F2048906B5056F042B;
defparam prom_inst_0.INIT_RAM_19 = 256'h0A91094B0B770F0E0EE809DD04D104A508330A5208FB07A309BF0D480D150800;
defparam prom_inst_0.INIT_RAM_1A = 256'h0FD50B050631063C09FF0C520B2C0A040C4D10000FF50B05061105FD09A10BD5;
defparam prom_inst_0.INIT_RAM_1B = 256'h077109F108FB08040A810E690E9509DD0524054A09290B990A9109870BEF0FC1;
defparam prom_inst_0.INIT_RAM_1C = 256'h06D70AB60ADC0623016B0197057F07FC0705060F088F0C7C0CAF080003510384;
defparam prom_inst_0.INIT_RAM_1D = 256'h000B000003B305FC04D403AE060109C409CF04FB002B003F04110679056F0467;
defparam prom_inst_0.INIT_RAM_1E = 256'h070505AE07CD0B5B0B2F0623011800F2048906B5056F042B065F0A0309EF04FB;
defparam prom_inst_0.INIT_RAM_1F = 256'h0EE809DD04D104A508330A5208FB07A309BF0D480D15080002EB02B80641085D;
defparam prom_inst_0.INIT_RAM_20 = 256'h09FF0C520B2C0A040C4D10000FF50B05061105FD09A10BD50A91094B0B770F0E;
defparam prom_inst_0.INIT_RAM_21 = 256'h0A810E690E9509DD0524054A09290B990A9109870BEF0FC10FD50B050631063C;
defparam prom_inst_0.INIT_RAM_22 = 256'h016B0197057F07FC0705060F088F0C7C0CAF080003510384077109F108FB0804;
defparam prom_inst_0.INIT_RAM_23 = 256'h04D403AE060109C409CF04FB002B003F04110679056F046706D70AB60ADC0623;
defparam prom_inst_0.INIT_RAM_24 = 256'h0B2F0623011800F2048906B5056F042B065F0A0309EF04FB000B000003B305FC;
defparam prom_inst_0.INIT_RAM_25 = 256'h08330A5208FB07A309BF0D480D15080002EB02B80641085D070505AE07CD0B5B;
defparam prom_inst_0.INIT_RAM_26 = 256'h0C4D10000FF50B05061105FD09A10BD50A91094B0B770F0E0EE809DD04D104A5;
defparam prom_inst_0.INIT_RAM_27 = 256'h0524054A09290B990A9109870BEF0FC10FD50B050631063C09FF0C520B2C0A04;
defparam prom_inst_0.INIT_RAM_28 = 256'h0705060F088F0C7C0CAF080003510384077109F108FB08040A810E690E9509DD;
defparam prom_inst_0.INIT_RAM_29 = 256'h09CF04FB002B003F04110679056F046706D70AB60ADC0623016B0197057F07FC;
defparam prom_inst_0.INIT_RAM_2A = 256'h048906B5056F042B065F0A0309EF04FB000B000003B305FC04D403AE060109C4;
defparam prom_inst_0.INIT_RAM_2B = 256'h09BF0D480D15080002EB02B80641085D070505AE07CD0B5B0B2F0623011800F2;
defparam prom_inst_0.INIT_RAM_2C = 256'h061105FD09A10BD50A91094B0B770F0E0EE809DD04D104A508330A5208FB07A3;
defparam prom_inst_0.INIT_RAM_2D = 256'h0A9109870BEF0FC10FD50B050631063C09FF0C520B2C0A040C4D10000FF50B05;
defparam prom_inst_0.INIT_RAM_2E = 256'h0CAF080003510384077109F108FB08040A810E690E9509DD0524054A09290B99;
defparam prom_inst_0.INIT_RAM_2F = 256'h04110679056F046706D70AB60ADC0623016B0197057F07FC0705060F088F0C7C;
defparam prom_inst_0.INIT_RAM_30 = 256'h065F0A0309EF04FB000B000003B305FC04D403AE060109C409CF04FB002B003F;
defparam prom_inst_0.INIT_RAM_31 = 256'h02EB02B80641085D070505AE07CD0B5B0B2F0623011800F2048906B5056F042B;
defparam prom_inst_0.INIT_RAM_32 = 256'h0A91094B0B770F0E0EE809DD04D104A508330A5208FB07A309BF0D480D150800;
defparam prom_inst_0.INIT_RAM_33 = 256'h0FD50B050631063C09FF0C520B2C0A040C4D10000FF50B05061105FD09A10BD5;
defparam prom_inst_0.INIT_RAM_34 = 256'h077109F108FB08040A810E690E9509DD0524054A09290B990A9109870BEF0FC1;
defparam prom_inst_0.INIT_RAM_35 = 256'h06D70AB60ADC0623016B0197057F07FC0705060F088F0C7C0CAF080003510384;
defparam prom_inst_0.INIT_RAM_36 = 256'h000B000003B305FC04D403AE060109C409CF04FB002B003F04110679056F0467;
defparam prom_inst_0.INIT_RAM_37 = 256'h070505AE07CD0B5B0B2F0623011800F2048906B5056F042B065F0A0309EF04FB;
defparam prom_inst_0.INIT_RAM_38 = 256'h0EE809DD04D104A508330A5208FB07A309BF0D480D15080002EB02B80641085D;
defparam prom_inst_0.INIT_RAM_39 = 256'h09FF0C520B2C0A040C4D10000FF50B05061105FD09A10BD50A91094B0B770F0E;
defparam prom_inst_0.INIT_RAM_3A = 256'h0A810E690E9509DD0524054A09290B990A9109870BEF0FC10FD50B050631063C;
defparam prom_inst_0.INIT_RAM_3B = 256'h016B0197057F07FC0705060F088F0C7C0CAF080003510384077109F108FB0804;
defparam prom_inst_0.INIT_RAM_3C = 256'h04D403AE060109C409CF04FB002B003F04110679056F046706D70AB60ADC0623;
defparam prom_inst_0.INIT_RAM_3D = 256'h0B2F0623011800F2048906B5056F042B065F0A0309EF04FB000B000003B305FC;
defparam prom_inst_0.INIT_RAM_3E = 256'h08330A5208FB07A309BF0D480D15080002EB02B80641085D070505AE07CD0B5B;
defparam prom_inst_0.INIT_RAM_3F = 256'h0C4D10000FF50B05061105FD09A10BD50A91094B0B770F0E0EE809DD04D104A5;

endmodule //fft_rom
