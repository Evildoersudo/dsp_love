//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.01 (64-bit)
//Part Number: GW5A-LV25UG324ES
//Device: GW5A-25
//Device Version: A
//Created Time: Sun Sep 22 20:41:30 2024

module fft_rom2 (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h08F908600B280F480F9E0B000647064B09E90C000A8D09030AD60E030D720800;
defparam prom_inst_0.INIT_RAM_01 = 256'h0B83062500D9007C03EC060C04D903C206370A310A8E062501CE025D06A8098A;
defparam prom_inst_0.INIT_RAM_02 = 256'h088B0B4E0A8D09B50C3310000FFB0B0005E9059408DD0AAA08F9074008F30C12;
defparam prom_inst_0.INIT_RAM_03 = 256'h07230A6C0A1705000005000003CD064B057304B207750BB10C43080003BD044F;
defparam prom_inst_0.INIT_RAM_04 = 256'h057205CF09C90C3E0B2709F40C140F840F2709DB047D03EE070D08C007070556;
defparam prom_inst_0.INIT_RAM_05 = 256'h05730400061709B509B90500006200B804D807A00707067609580DA30E3209DB;
defparam prom_inst_0.INIT_RAM_06 = 256'h0F9E0B000647064B09E90C000A8D09030AD60E030D720800028E01FD052A06FD;
defparam prom_inst_0.INIT_RAM_07 = 256'h03EC060C04D903C206370A310A8E062501CE025D06A8098A08F908600B280F48;
defparam prom_inst_0.INIT_RAM_08 = 256'h0C3310000FFB0B0005E9059408DD0AAA08F9074008F30C120B83062500D9007C;
defparam prom_inst_0.INIT_RAM_09 = 256'h0005000003CD064B057304B207750BB10C43080003BD044F088B0B4E0A8D09B5;
defparam prom_inst_0.INIT_RAM_0A = 256'h0B2709F40C140F840F2709DB047D03EE070D08C00707055607230A6C0A170500;
defparam prom_inst_0.INIT_RAM_0B = 256'h09B90500006200B804D807A00707067609580DA30E3209DB057205CF09C90C3E;
defparam prom_inst_0.INIT_RAM_0C = 256'h09E90C000A8D09030AD60E030D720800028E01FD052A06FD05730400061709B5;
defparam prom_inst_0.INIT_RAM_0D = 256'h06370A310A8E062501CE025D06A8098A08F908600B280F480F9E0B000647064B;
defparam prom_inst_0.INIT_RAM_0E = 256'h05E9059408DD0AAA08F9074008F30C120B83062500D9007C03EC060C04D903C2;
defparam prom_inst_0.INIT_RAM_0F = 256'h057304B207750BB10C43080003BD044F088B0B4E0A8D09B50C3310000FFB0B00;
defparam prom_inst_0.INIT_RAM_10 = 256'h0F2709DB047D03EE070D08C00707055607230A6C0A1705000005000003CD064B;
defparam prom_inst_0.INIT_RAM_11 = 256'h04D807A00707067609580DA30E3209DB057205CF09C90C3E0B2709F40C140F84;
defparam prom_inst_0.INIT_RAM_12 = 256'h0AD60E030D720800028E01FD052A06FD05730400061709B509B90500006200B8;
defparam prom_inst_0.INIT_RAM_13 = 256'h01CE025D06A8098A08F908600B280F480F9E0B000647064B09E90C000A8D0903;
defparam prom_inst_0.INIT_RAM_14 = 256'h08F9074008F30C120B83062500D9007C03EC060C04D903C206370A310A8E0625;
defparam prom_inst_0.INIT_RAM_15 = 256'h0C43080003BD044F088B0B4E0A8D09B50C3310000FFB0B0005E9059408DD0AAA;
defparam prom_inst_0.INIT_RAM_16 = 256'h070D08C00707055607230A6C0A1705000005000003CD064B057304B207750BB1;
defparam prom_inst_0.INIT_RAM_17 = 256'h09580DA30E3209DB057205CF09C90C3E0B2709F40C140F840F2709DB047D03EE;
defparam prom_inst_0.INIT_RAM_18 = 256'h028E01FD052A06FD05730400061709B509B90500006200B804D807A007070676;
defparam prom_inst_0.INIT_RAM_19 = 256'h08F908600B280F480F9E0B000647064B09E90C000A8D09030AD60E030D720800;
defparam prom_inst_0.INIT_RAM_1A = 256'h0B83062500D9007C03EC060C04D903C206370A310A8E062501CE025D06A8098A;
defparam prom_inst_0.INIT_RAM_1B = 256'h088B0B4E0A8D09B50C3310000FFB0B0005E9059408DD0AAA08F9074008F30C12;
defparam prom_inst_0.INIT_RAM_1C = 256'h07230A6C0A1705000005000003CD064B057304B207750BB10C43080003BD044F;
defparam prom_inst_0.INIT_RAM_1D = 256'h057205CF09C90C3E0B2709F40C140F840F2709DB047D03EE070D08C007070556;
defparam prom_inst_0.INIT_RAM_1E = 256'h05730400061709B509B90500006200B804D807A00707067609580DA30E3209DB;
defparam prom_inst_0.INIT_RAM_1F = 256'h0F9E0B000647064B09E90C000A8D09030AD60E030D720800028E01FD052A06FD;
defparam prom_inst_0.INIT_RAM_20 = 256'h03EC060C04D903C206370A310A8E062501CE025D06A8098A08F908600B280F48;
defparam prom_inst_0.INIT_RAM_21 = 256'h0C3310000FFB0B0005E9059408DD0AAA08F9074008F30C120B83062500D9007C;
defparam prom_inst_0.INIT_RAM_22 = 256'h0005000003CD064B057304B207750BB10C43080003BD044F088B0B4E0A8D09B5;
defparam prom_inst_0.INIT_RAM_23 = 256'h0B2709F40C140F840F2709DB047D03EE070D08C00707055607230A6C0A170500;
defparam prom_inst_0.INIT_RAM_24 = 256'h09B90500006200B804D807A00707067609580DA30E3209DB057205CF09C90C3E;
defparam prom_inst_0.INIT_RAM_25 = 256'h09E90C000A8D09030AD60E030D720800028E01FD052A06FD05730400061709B5;
defparam prom_inst_0.INIT_RAM_26 = 256'h06370A310A8E062501CE025D06A8098A08F908600B280F480F9E0B000647064B;
defparam prom_inst_0.INIT_RAM_27 = 256'h05E9059408DD0AAA08F9074008F30C120B83062500D9007C03EC060C04D903C2;
defparam prom_inst_0.INIT_RAM_28 = 256'h057304B207750BB10C43080003BD044F088B0B4E0A8D09B50C3310000FFB0B00;
defparam prom_inst_0.INIT_RAM_29 = 256'h0F2709DB047D03EE070D08C00707055607230A6C0A1705000005000003CD064B;
defparam prom_inst_0.INIT_RAM_2A = 256'h04D807A00707067609580DA30E3209DB057205CF09C90C3E0B2709F40C140F84;
defparam prom_inst_0.INIT_RAM_2B = 256'h0AD60E030D720800028E01FD052A06FD05730400061709B509B90500006200B8;
defparam prom_inst_0.INIT_RAM_2C = 256'h01CE025D06A8098A08F908600B280F480F9E0B000647064B09E90C000A8D0903;
defparam prom_inst_0.INIT_RAM_2D = 256'h08F9074008F30C120B83062500D9007C03EC060C04D903C206370A310A8E0625;
defparam prom_inst_0.INIT_RAM_2E = 256'h0C43080003BD044F088B0B4E0A8D09B50C3310000FFB0B0005E9059408DD0AAA;
defparam prom_inst_0.INIT_RAM_2F = 256'h070D08C00707055607230A6C0A1705000005000003CD064B057304B207750BB1;
defparam prom_inst_0.INIT_RAM_30 = 256'h09580DA30E3209DB057205CF09C90C3E0B2709F40C140F840F2709DB047D03EE;
defparam prom_inst_0.INIT_RAM_31 = 256'h028E01FD052A06FD05730400061709B509B90500006200B804D807A007070676;
defparam prom_inst_0.INIT_RAM_32 = 256'h08F908600B280F480F9E0B000647064B09E90C000A8D09030AD60E030D720800;
defparam prom_inst_0.INIT_RAM_33 = 256'h0B83062500D9007C03EC060C04D903C206370A310A8E062501CE025D06A8098A;
defparam prom_inst_0.INIT_RAM_34 = 256'h088B0B4E0A8D09B50C3310000FFB0B0005E9059408DD0AAA08F9074008F30C12;
defparam prom_inst_0.INIT_RAM_35 = 256'h07230A6C0A1705000005000003CD064B057304B207750BB10C43080003BD044F;
defparam prom_inst_0.INIT_RAM_36 = 256'h057205CF09C90C3E0B2709F40C140F840F2709DB047D03EE070D08C007070556;
defparam prom_inst_0.INIT_RAM_37 = 256'h05730400061709B509B90500006200B804D807A00707067609580DA30E3209DB;
defparam prom_inst_0.INIT_RAM_38 = 256'h0F9E0B000647064B09E90C000A8D09030AD60E030D720800028E01FD052A06FD;
defparam prom_inst_0.INIT_RAM_39 = 256'h03EC060C04D903C206370A310A8E062501CE025D06A8098A08F908600B280F48;
defparam prom_inst_0.INIT_RAM_3A = 256'h0C3310000FFB0B0005E9059408DD0AAA08F9074008F30C120B83062500D9007C;
defparam prom_inst_0.INIT_RAM_3B = 256'h0005000003CD064B057304B207750BB10C43080003BD044F088B0B4E0A8D09B5;
defparam prom_inst_0.INIT_RAM_3C = 256'h0B2709F40C140F840F2709DB047D03EE070D08C00707055607230A6C0A170500;
defparam prom_inst_0.INIT_RAM_3D = 256'h09B90500006200B804D807A00707067609580DA30E3209DB057205CF09C90C3E;
defparam prom_inst_0.INIT_RAM_3E = 256'h09E90C000A8D09030AD60E030D720800028E01FD052A06FD05730400061709B5;
defparam prom_inst_0.INIT_RAM_3F = 256'h06370A310A8E062501CE025D06A8098A08F908600B280F480F9E0B000647064B;

endmodule //fft_rom2
